
module unsaved (
	);	

endmodule
