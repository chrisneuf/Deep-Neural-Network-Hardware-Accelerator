module tb_dnn_bonus();
endmodule: tb_dnn_bonus
